class generator;

    transaction tr;
    mailbox #(transaction) mbx;
    event done;
    int count = 0;
    event drvnext;
    event sconext;

    function new(mailbox #(transaction) mbx);
        this.mbx = mbx;
        tr = new();
    endfunction

    task run();
        repeat(count) begin
            assert(tr.randomize) else $error("[GEN] Randomization Failed");
            mbx.put(tr.copy);
            $display("[GEN]: Oper : %0s Din : %0d", tr.oper.name(), tr.dintx);
            @(drvnext);
            @(sconext);
        end
        -> done;
    endtask

endclass
